`include "Rsa256Core.sv"
