`include "Rsa256Core.sv"
`include "Rsa256Wrapper.sv"
